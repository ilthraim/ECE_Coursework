module rcvr_top(

    );
endmodule
