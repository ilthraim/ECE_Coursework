module xmit_controller(
    input logic clk, rst, xvalid, cardet, mx_rdy, xsend, ack_needed, ack_recieved, [7:0] mac,
    output logic xrdy, mx_valid, [7:0] xerrcnt);
    
    
    
endmodule
