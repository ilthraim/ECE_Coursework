module FinalProjectTop(
    input logic clk, rst, uart_in, rxd, [7:0] mac, [1:0] f_type, [1:0] dest,
    output logic uart_out, txen, txd, cfgdat, dp_n, [7:0] an_n, [6:0] segs_n);
    
    
    
endmodule
