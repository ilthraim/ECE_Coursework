module xmit_top #(parameter BIT_RATE = 50000) (
    input logic clk, rst, cardet, ACK_recieved, ACK_needed, [7:0] mac, ack_addr, [1:0] dest_addr, ftype, uart_in,
    output logic [7:0] xerrcnt);

    

endmodule